`ifndef APB_ENV
`define APB_ENV
class apb_env extends uvm_env;
  `uvm_component_utils(apb_env)
  apb_agent agt;
  apb_scoreboard scb;
  function new(string name = "apb_env", uvm_component parent);
    super.new(name,parent);
  endfunction
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    agt = apb_agent::type_id::create("agt", this);
    scb = apb_scoreboard::type_id::create("scb", this);
  endfunction
  function void connect_phase(uvm_phase phase);
    agt.mon.mon_ap.connect(scb.sb_imp);
  endfunction
endclass
`endif
